`timescale 1ns / 1ps 
// `include "clogb2.v" // vivado can't find this for some reason
//////////////////////////////////////////////////////////////////////////////////
// Copyright (c) Gyorgy Wyatt Muntean 2017
// Create Date: 02/25/2017 12:04:27 PM
// Module Name: dotProduct_testbench
// Project Name: Matrix Multiply
// Target Devices: ZYNQ702
// Description: 
//      This module serves as a testbench for the dotProduct module.
//
//////////////////////////////////////////////////////////////////////////////////

module dotProduct_testbench2();
    localparam DIM = 22;
    localparam A_DATA_WIDTH = 32;
    localparam B_DATA_WIDTH = 32;
    localparam EXTRA_ADD_WIDTH =  5;    //`CLOG2(DIM); // this isnt working for now...
    localparam RES_WIDTH = A_DATA_WIDTH + B_DATA_WIDTH + EXTRA_ADD_WIDTH;
    
    reg Clock;
    reg start;
    reg [(A_DATA_WIDTH*DIM)-1:0] A;
    reg [(B_DATA_WIDTH*DIM)-1:0] B;
    wire [RES_WIDTH-1:0] DotProduct;
    wire readEn;
    
    // Set up the clock.
    parameter CLOCK_PERIOD=10;
    initial Clock=1;
    always begin
        #(CLOCK_PERIOD/2);
        Clock = ~Clock;
    end
    
    // unit under test
    dotProduct #(DIM, A_DATA_WIDTH, B_DATA_WIDTH, RES_WIDTH) uut(.Clock(Clock), .start(start), .A(A), .B(B), .DotProduct(DotProduct), .readEn(readEn) );    
    
    // Try silly input case
    initial begin  
			// Initialize inputs
			A = 0;
			B = 0;

			@(posedge Clock);
			@(posedge Clock);
			@(posedge Clock);
			@(posedge Clock);
			@(posedge Clock);
			@(posedge Clock);

			A = 704'b11011000000001110010101111001100101011010011000110001001100001111101011101110000110111000111000101010000010000010010100010101011101101000000100001011101000011111110111100110100111101011110000111001000110000001110100000000111111110000111111010110000000111111011110011001001000001000010010110001101111101110101010011101010110010011011110100010101011110000011001010011101110101100000101110110010100010110000000011110010001101101111111000101100111101010110111010100101001110110110111001011111010001010100000110100101010100001011110100011111110111101010010100000100001000111000011011010101001101111100010110010111111011101000001001110001101101011101110010111010010000110100001100101000100001101110001001000000;
			B = 704'b01000010000001100100000100111010011011101100011010100101110100101111101010100101110111010110010011101010101001110011100111001010111110111101101001001100010110100001000100100010100110110001110011011111000000011001011000110010100010110011011100001000000010001001111101101101000100100011100100001101010010010110100000001001001100011000110100111100001100011010000000100010111000010001101110000101000101011001001001001101101001101110010100010001111101010010110100101101110001010010011100000101000001101111000110101101100001100100001011100001010100011011111110111111111010101010001010101101000010101001100010110111011001010100110101101101100001000110010110110000100100110000010011011111100111100101111010000101;
			// Expected result = 129094160280529530105
			start = 1; @(posedge Clock)
			start = 0; @(posedge Clock)
			A = 704'b10011011100011100100011110111001111111010000110100000111111110000101011100100100001111000000011011101010010111001111101011001010011110001000010111000111101100111010011101111101110010111010010111101101111010011100000010111011101110110010010110000001110111101011101111001111101111111101000101011010100011110101100010000000001100110111000101001001000101100011111110111110111001011110000111000110010000101111110000010110001000111011101001011101011111110010010101000010101011101101000100110111111000001100000110010101011001101100100001110101110110111001000100011111100001010011001011001011011000100000001110101101101001111000111110010010111101100100000010001100110111101001011010111110001010100110101000011110;
			B = 704'b01110010011001100110110101101000011000011011000110110101010011111000010000101011010110101101101100001010101110100010111011101110011111110111011010011100100110100011010111101101000001000110101000110000010011111110110000100010010001010001010000101011100011100001001011110101010110100111111100110100101111010101100011111110111110010011010011101100010000011101110000101001010000111101000110111100001110110000111100110011110010001001001111111101011101101010011110111111000100010111011000110010011111110100101010111001110011111000100010000101110001111001011000100111011001100100111000000100001110001010000011111110000111011010111101011101000100010010101110000010000010100101110011001100100110111100111110011010;
			// Expected result = 80159935725743712742
			start = 1; @(posedge Clock)
			start = 0; @(posedge Clock)
			A = 704'b01111110110100110001001111111110010011001100000101111011011100011111011000010100101011100101101111100110110101100001100111100101101000110111110100101010011000000111100111101110000000100101001101110110011100000011101110111101101110111110010100011000000100100010000011011011100011001101001100001011001101100110001010001111010101011000100000111101100000111100000011000110010111011110010011010001010111000110110000111101011110100001000110100010100000101101000010100101001100010000011010111010001111001000011001011100011001110111101100111100101100110110000011100110000000011011011000111110001000001000100000001011111110000101001011000111111010110110100101110101110001011010011010010010010011010111101010101010;
			B = 704'b00101111010100000101000101000000001100100110011111001100101000000010110011110011111110101010001011000001010111011001110001010001000100110001101001000000000110000100101010001001001001011001101010011011110000111110010001111001011110100001000001000010100110111101001000011110100001000110110000101111111100101111000110000011101110100011100111100110100101110101010101010011001100001111011000000000101111101100010000001011001100100101100111111111110010010010110010001010010011110100000000101001100110101000000101011101010101010000110101110110100111100110101000110100100101000111110100010011000000001011010110110111101110010000001000010100011110000101000111100101100101010001010110100010001110001001011000001011;
			// Expected result = 79068974242824022472
			start = 1; @(posedge Clock)
			start = 0; @(posedge Clock)
			A = 704'b10001100110010011111101011101001001001111010111111111011010111100111001111010000001111010010101100100000011100111110010100000111110110110000110110001111011111010100111100101010001101100111101000011001111110011101010001000011110100001010001001101111010110111001101101001111111110001011110010101000111001011111010111000110001111001100001000001100001100011000000110111110010100010111010101001010010010101101100111010100111001010001000001100001001101001110010000110111000001101100110100100001100110011000011011000110001101001010100110000110001010100000100111100100100100100110100000101000000011011011010000100111001111111101101010001111100001100101110111110000010110000001110111100011100110101010100011111000;
			B = 704'b01100110101110100000010110011001011101000001100101011110001101001110000111101011010011101001001010010100110001101100011001111101101110110011000110101101101010101111111100011001000101011111011111111110110000110010011001111111000010101010110001010000110110110000110000000010011000101111111100010101001000111001010001110101010101011010010000000100101111111111000001111101100011101010100110011110100101110100110110100110101110111000011110001000011100011101000100111100110010001100000111101111010010111100011010011001111100110011101111100010011111010100010000001010110111000110100011011110111001011100100111000101001101001011000011110001011010110000000101001011101010001110101011010100111011100101101001010010;
			// Expected result = 97626475732690395310
			start = 1; @(posedge Clock)
			start = 0; @(posedge Clock)
			A = 704'b11011111110101100000000001011100100111010110100111110001101010000100000001111011000110010101010001100100100000100010011001110111000011110000010101111111000010111001111011011001111111110010000110111110010101001101101101001010100000010110111010101010110000000110001101011010110101100001001000000011110101101011101001000101101010011111010110011101011000110010110100011001111000100100101011100100100111011111011011101010000100001011011101111000111111010011110111110101110010100100110111101011101111010000100111010001100101110011111101011101111010101100101100111011010100101011101100111101111111101100100100001011110001011110001101111110111100001110110000000001001111111001001111110111010110100001111000110111;
			B = 704'b10111100111100011111101111001111001010111101010101100000100110110110111001001010111101010001101110000011000100110000101011001100001111111100010101110001110111100011111110110010100000001101110000101010010110001111101111101011011111111100010001000010101001110111000010100110000011000010101010011101100001110101100101010001001111001100101100010111001000110111011001001000110001111010011011011001100011011011100101110011110001011101110100100001100110011010010011010010101000100001010011111101011110011011101001001011010101000110101010101011000111100001000000011101101101010011111011001011111110101001100111100101101101101111101100111111111101100100100101101011011110110000110000111010110101111101011010110110;
			// Expected result = 99193988133750016235
			start = 1; @(posedge Clock)
			start = 0; @(posedge Clock)
			A = 704'b10011110101011100101101100111100010111100111001110110110011111110001001111111111111110011101101000111010110100101110001010101100111010101110001001011110000111100110011001100011001010111110011111001011011010110001101001101001010101101111001010000010011111001011100100001100111000000000011010100001001010101111001001100001010101100100111010001000101111000010011010001000110111000000101101011110010010111011111101100011000111111010010000110110010110000101101000010101011001110101111001111001110100111000101111111101111011110111001011000010001001010000010110000100100000000010101010001100010111001010100000101100110011010001011001101010110110011110101011010010001001000000000101000010010011011100100101101101;
			B = 704'b00101001100010001101100001111000101110101010100010000000011110011101010011111111110111001000011010111011110110000101110101011001111110010100000011010100011001110011111110101010001000000010101100101100000111000101101000001000110101010000000110111111110000100111000000000001100010101010110000100000000010001101100000000101110011000100000101111100001010011001000100110100100100101101001001100000010010110011000100111010001000111010010100001100110011010000011111011101110110101100101010101110101101000100100001111110001101111101101000100111110001000110111101011111010000000101000101011010111000111100110100111101101001101010010001110110101010000010100001001001011000001001111110100111100110111001011111101100;
			// Expected result = 83006198284222388338
			start = 1; @(posedge Clock)
			start = 0; @(posedge Clock)
			A = 704'b00000100100110111001000001011110100100111101110110110000001111011000110000011000111101001010010111100000101110100111110100111010010010100110100101010011110011110010111111011100001000101010011101000010011001000100111100000101011111010100111111111010001000000010001101100100000010011111010110001010001000111010010110110010010110010111100110101000001101101011100110011010001100111101011011000110001100101011001010110100110110000111011010000110111100001001100110111111010000011000101000010110111001101110110111101111010010001011110010100010111101111110100100000111001011111101111100100001001111111110100111010011111010100111011110100110101001011110101001000110011111101001101100101111110110110101110010010010;
			B = 704'b11000001101100110101010111110010100010000100101000110011001010010011011010100111011101001010100001110110000010001101011010010010000101010001100010011111011011001111001111000101111010010011010101110110000001110100011010101110011010000100011111000010001011010100111010001110110111011110101100010001001010001100100100111101001110011000010110101100101001110100000001101010100000100111010010111101110100101101010101010011100011001101101010100010100011011111010010001011110111011100011001010011000000101000101010111100001101101000100011000111100100110110111010000110001100110111100000100010001001101100000001111001110110011111001011010010001100011001000010111011011011001101000001100100001110100011110101011011;
			// Expected result = 95672266352123932092
			start = 1; @(posedge Clock)
			start = 0; @(posedge Clock)
			A = 704'b01110110111111100011100111000010110101110010011000001110011000100111001111010001111100011000100101101100111000101100100010110101010110001001111110011000110010100011111100100100101010000111100001000000011000001111001001100011110000100100100001100011100100000111111101010001100100111000010011001000111001000000011111111110110001001010011110111111111101010101010100110100011001011001010101000111011110111010000100011011010000010100010001100110011000010011100010011100111011111000110110011010100011100001110010001111001110111111110100100001010001010101000101001001100000111101111110101011101001001100010110001100011100000111111111000110111101110100001101000110100001101001010001011011101000011110100001101011;
			B = 704'b10100010111101111011011001001010111001100010000010100101111110011010100110111010000001101001111100010001011110100110010101010011110010100100000001010100101010001001101101101100001111010010100101111000110101001111000011011011000011100000010011110011010101100000011010010010110010011101011100010011100010000111101001100101101100010101011101100000000101111001100010100101000100010101110101111111000110001100100111110111101000111111111101101011000110010110000100100110011001001100011110101011110100000000011100011001101000011011100001110011010011001011000010000011111110001000101011111111101101000011011010110111010101110111100000011111100111100111111000100101000011001011001110000010010010110111000000100010;
			// Expected result = 93279828370341815357
			start = 1; @(posedge Clock)
			start = 0; @(posedge Clock)
			A = 704'b00100110101101111011001100001010011000001010111000100111101110101111000011011011010001101011001111010001010010001001101100000010010010111000011110010000111110110110110110010100000100011000111010011111001010100000010000111000001000111010000100101101100111001101001101111000010100001111101011000010101100110110010011100010110010111111000010010010001101001111001111111000011110111000101101110011111000001000000000011100000010011111100000100000011011010100101101100000000000000001010111001001110001111100101011000001110000000101101001100110101100101000010100110100010000011100000010000001000000011010001100111000010011110001110100001100100000000011000100010001001100100111111111000011110111000111011010111001;
			B = 704'b01110101110011001110001011001100011011001010001000011001101010011010001011010011110111011101001100001111110001000001110100001110000110010100101010111110011010010011100000000010100001111001101011101010111011111000001110110100110111110001001001100010000010010101010111011001111101011111011101100111110111111011111111111010100100101100001100011111111001101001000110110001111110111110111001010100110100100100001101010111101111100110010111111101110101100110001110111010101100101011101000011101100100001111011110111101111010100010100110011100010011111010010100010000100100001110110100000011111110010000011111100110000100011011011110100101101001000100001110111001010101101000000111101101000000111101011111001101;
			// Expected result = 100971865087261433601
			start = 1; @(posedge Clock)
			start = 0; @(posedge Clock)
			A = 704'b10110111100111111010111100011000011100011100110110000011001000100111101000100110110111110100011100100000111110011111100000111100000110010010101000110000101101011110001110110000000111001011100100000011110011101000101011001101100111011000101111001111010101111011101101101110000000111100101110110000111001111111100010000010101010110101101010110100011101101010011011010000000000111001010110110011110010100011111100011111011001111011001101000000000111110011110110011110111010000110001010110111010101101110011001011100101101010010110011011110001011110110001101000110110000111000111111110010000011100000110011101011000101111010101000000110111011101001010001110101110001111110100001100100001011100111110000001110;
			B = 704'b10000110101110110000011110110010110011010010010111010101101011001001010000001101100111011000110100110111111100110000011001110001010100001111010011101110001111101011101011000101111101111001001110011011011010000000010001111101101101111110111001110010011001001101011101111001000010101001111001101101100100001011001000011011100000100010010000010011011001011010000110011101001011101001000010010110000100001011000100100011101110011101111011001010101011100001011111100001001001110101010110011010110111111100010100110010010111111001110100110101110001110110011110111000011101011110000111000011010111000001000010001101101111001010001110110100010001100000101010111111111001001111011111100010110101111011101000000000;
			// Expected result = 121313163178808512007
			start = 1; @(posedge Clock)
			start = 0; @(posedge Clock)
			#100;
		end 
endmodule
