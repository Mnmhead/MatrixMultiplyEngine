`timescale 1ns / 1ps 
// `include "clogb2.v" // vivado can't find this for some reason
//////////////////////////////////////////////////////////////////////////////////
// Copyright (c) Gyorgy Wyatt Muntean 2017
// Create Date: 02/25/2017 12:04:27 PM
// Module Name: dotProduct_testbench
// Project Name: Matrix Multiply
// Target Devices: ZYNQ702
// Description: 
//      This module serves as a testbench for the dotProduct module.
//
//////////////////////////////////////////////////////////////////////////////////

module dotProduct_testbench();
    localparam DIM = 10;
    localparam A_DATA_WIDTH = 16;
    localparam B_DATA_WIDTH = 16;
    localparam EXTRA_ADD_WIDTH =  4;    //`CLOG2(DIM); // this isnt working for now...
    localparam RES_WIDTH = A_DATA_WIDTH + B_DATA_WIDTH + EXTRA_ADD_WIDTH;
    
    reg Clock;
    reg [(A_DATA_WIDTH*DIM)-1:0] A;
    reg [(B_DATA_WIDTH*DIM)-1:0] B;
    wire [RES_WIDTH-1:0] DotProduct;
    
    // Set up the clock.
    parameter CLOCK_PERIOD=10;
    initial Clock=1;
    always begin
        #(CLOCK_PERIOD/2);
        Clock = ~Clock;
    end
    
    // unit under test
    dotProduct #(DIM, A_DATA_WIDTH, B_DATA_WIDTH) uut(.Clock(Clock), .A(A), .B(B), .DotProduct(DotProduct));    
    
    // Try silly input case
    initial begin  
        // Initialize inputs
        A = 0;
        B = 0;
        
        // pause for 100 ns
        #100;  
        
        A = 160'b0000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000;
        B = 160'b0000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000;
        // Expected result = 640
        @(posedge Clock);
        @(posedge Clock);
        A = 160'b1001011100100101101101010100000101000001111001110001101101001011011100111100000111001010000000000111000101100111010000110100000111111110110001011111011101111000;
        B = 160'b1010011111010001010000111101011011001111111011001100001010010110101101000100000010110001001100010111110110110001010100101101011101010001000001101101110101011110;
        // Expected result = 13669466157
        @(posedge Clock)
        @(posedge Clock)
        A = 160'b1111001010000001110010100000000001110001011001000000110011100100001101111110110101000001110000010001000101000101010000100110100100111110100011101111001100111000;
        B = 160'b0010000011111111000111000011000010001010100110011000001011101000111011001001111001100001111110001110100111000110111110100100000000001110100010001100111001101001;
        // Expected result = 8030888999
        @(posedge Clock)
        @(posedge Clock)
        A = 160'b1100101001000010110010001111111000001010111101001110011011001011100001101101111001101101100111100111101100101100101011101111111111111111111101000000110110101111;
        B = 160'b0111100001010001101110110000110101101010010001000000111100101000110100101000011011011001010101111100100001010101100001011011100000011010001111111001110100011111;
        // Expected result = 11518131799
        @(posedge Clock)
        @(posedge Clock)
        A = 160'b0101100011100011111100100100101001010011011000001001101110011001010001111110011111010101111111100000001111111011111001001010111100100101111110000011100101111001;
        B = 160'b1010001011101100000100011101001111111110000001000010101000001110101000110000101000110011010011001000010110000111100110010010111001101110101011101111110000110000;
        // Expected result = 8092373917
        @(posedge Clock)
        @(posedge Clock)
        A = 160'b0011011010011111111110011011111100001001100000000001010100010011001100101000001101100100010111111010101110111111110000101000111101001111110110100001110101100110;
        B = 160'b0100001000000111100001000110000001001001011000011011101000010000100101111110000100100100100011011101110010101101101011000000010111101011000111010101010110101000;
        // Expected result = 9521434271
        @(posedge Clock)
        @(posedge Clock)
        A = 160'b0111001010100110100101100101010100101101111001000011010111000111001010100010011111100100111000101010111010101010001000010001111001110111011100011001100110010000;
        B = 160'b0101111100001111000010000001100010111110111101010111010101000111100100100110111100100110010110011001000010101100001000111101110101101010110010011011011110010010;
        // Expected result = 7178516105
        @(posedge Clock)
        @(posedge Clock)
        A = 160'b1000011000000000100011110000101100011010101011110001001111111101111000111110010111101111000110000100100110110111001100010111110101011110101001111010011111100010;
        B = 160'b0001011000111100111100011100001000111100001110011100000100100010011010110101000110100100010100111010010100001100010001010111001111011000001100001010011000101011;
        // Expected result = 11189416997
        @(posedge Clock)
        @(posedge Clock)
        A = 160'b0000101000101101011001111100110111101011101110000001111010110010110001010001001011000000100110010101100110101111110100011000011100010001100100111100101000000001;
        B = 160'b0110011111101001001010100010001011100111101100110100001101011111110100110100010000011101001110010011000110100011100111110001011000111101001101101001101011000010;
        // Expected result = 11763638665
        
        #100;
    end 
endmodule
